module chess

pub const pawn_attacks = [
	[Bitboard(0)],
	[Bitboard(0x200), 0x500, 0xa00, 0x1400, 0x2800, 0x5000, 0xa000, 0x4000, 0x20000, 0x50000, 0xa0000,
		0x140000, 0x280000, 0x500000, 0xa00000, 0x400000, 0x2000000, 0x5000000, 0xa000000, 0x14000000,
		0x28000000, 0x50000000, 0xa0000000, 0x40000000, 0x200000000, 0x500000000, 0xa00000000,
		0x1400000000, 0x2800000000, 0x5000000000, 0xa000000000, 0x4000000000, 0x20000000000,
		0x50000000000, 0xa0000000000, 0x140000000000, 0x280000000000, 0x500000000000, 0xa00000000000,
		0x400000000000, 0x2000000000000, 0x5000000000000, 0xa000000000000, 0x14000000000000,
		0x28000000000000, 0x50000000000000, 0xa0000000000000, 0x40000000000000, 0x200000000000000,
		0x500000000000000, 0xa00000000000000, 0x1400000000000000, 0x2800000000000000,
		0x5000000000000000, 0xa000000000000000, 0x4000000000000000, 0x0, 0x0, 0x0, 0x0, 0x0, 0x0,
		0x0, 0x0],
	[Bitboard(0x0), 0x0, 0x0, 0x0, 0x0, 0x0, 0x0, 0x0, 0x2, 0x5, 0xa, 0x14, 0x28, 0x50, 0xa0, 0x40,
		0x200, 0x500, 0xa00, 0x1400, 0x2800, 0x5000, 0xa000, 0x4000, 0x20000, 0x50000, 0xa0000,
		0x140000, 0x280000, 0x500000, 0xa00000, 0x400000, 0x2000000, 0x5000000, 0xa000000, 0x14000000,
		0x28000000, 0x50000000, 0xa0000000, 0x40000000, 0x200000000, 0x500000000, 0xa00000000,
		0x1400000000, 0x2800000000, 0x5000000000, 0xa000000000, 0x4000000000, 0x20000000000,
		0x50000000000, 0xa0000000000, 0x140000000000, 0x280000000000, 0x500000000000, 0xa00000000000,
		0x400000000000, 0x2000000000000, 0x5000000000000, 0xa000000000000, 0x14000000000000,
		0x28000000000000, 0x50000000000000, 0xa0000000000000, 0x40000000000000],
]

pub const knight_attacks = [
	Bitboard(0x20400),
	0x50800,
	0xa1100,
	0x142200,
	0x284400,
	0x508800,
	0xa01000,
	0x402000,
	0x2040004,
	0x5080008,
	0xa110011,
	0x14220022,
	0x28440044,
	0x50880088,
	0xa0100010,
	0x40200020,
	0x204000402,
	0x508000805,
	0xa1100110a,
	0x1422002214,
	0x2844004428,
	0x5088008850,
	0xa0100010a0,
	0x4020002040,
	0x20400040200,
	0x50800080500,
	0xa1100110a00,
	0x142200221400,
	0x284400442800,
	0x508800885000,
	0xa0100010a000,
	0x402000204000,
	0x2040004020000,
	0x5080008050000,
	0xa1100110a0000,
	0x14220022140000,
	0x28440044280000,
	0x50880088500000,
	0xa0100010a00000,
	0x40200020400000,
	0x204000402000000,
	0x508000805000000,
	0xa1100110a000000,
	0x1422002214000000,
	0x2844004428000000,
	0x5088008850000000,
	0xa0100010a0000000,
	0x4020002040000000,
	0x400040200000000,
	0x800080500000000,
	0x1100110a00000000,
	0x2200221400000000,
	0x4400442800000000,
	0x8800885000000000,
	0x100010a000000000,
	0x2000204000000000,
	0x4020000000000,
	0x8050000000000,
	0x110a0000000000,
	0x22140000000000,
	0x44280000000000,
	0x88500000000000,
	0x10a00000000000,
	0x20400000000000,
]

pub const king_attacks = [
	Bitboard(0x302),
	0x705,
	0xe0a,
	0x1c14,
	0x3828,
	0x7050,
	0xe0a0,
	0xc040,
	0x30203,
	0x70507,
	0xe0a0e,
	0x1c141c,
	0x382838,
	0x705070,
	0xe0a0e0,
	0xc040c0,
	0x3020300,
	0x7050700,
	0xe0a0e00,
	0x1c141c00,
	0x38283800,
	0x70507000,
	0xe0a0e000,
	0xc040c000,
	0x302030000,
	0x705070000,
	0xe0a0e0000,
	0x1c141c0000,
	0x3828380000,
	0x7050700000,
	0xe0a0e00000,
	0xc040c00000,
	0x30203000000,
	0x70507000000,
	0xe0a0e000000,
	0x1c141c000000,
	0x382838000000,
	0x705070000000,
	0xe0a0e0000000,
	0xc040c0000000,
	0x3020300000000,
	0x7050700000000,
	0xe0a0e00000000,
	0x1c141c00000000,
	0x38283800000000,
	0x70507000000000,
	0xe0a0e000000000,
	0xc040c000000000,
	0x302030000000000,
	0x705070000000000,
	0xe0a0e0000000000,
	0x1c141c0000000000,
	0x3828380000000000,
	0x7050700000000000,
	0xe0a0e00000000000,
	0xc040c00000000000,
	0x203000000000000,
	0x507000000000000,
	0xa0e000000000000,
	0x141c000000000000,
	0x2838000000000000,
	0x5070000000000000,
	0xa0e0000000000000,
	0x40c0000000000000,
]

pub const ray_attacks = [
	[
		Bitboard(0x0),
		0x0,
		0x2,
		0x6,
		0xE,
		0x1E,
		0x3E,
		0x7E,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x100,
		0x0,
		0x200,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x10100,
		0x0,
		0x0,
		0x40200,
		0x0,
		0x0,
		0x0,
		0x0,
		0x1010100,
		0x0,
		0x0,
		0x0,
		0x8040200,
		0x0,
		0x0,
		0x0,
		0x101010100,
		0x0,
		0x0,
		0x0,
		0x0,
		0x1008040200,
		0x0,
		0x0,
		0x10101010100,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x201008040200,
		0x0,
		0x1010101010100,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40201008040200,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x4,
		0xC,
		0x1C,
		0x3C,
		0x7C,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x200,
		0x0,
		0x400,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20200,
		0x0,
		0x0,
		0x80400,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2020200,
		0x0,
		0x0,
		0x0,
		0x10080400,
		0x0,
		0x0,
		0x0,
		0x202020200,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2010080400,
		0x0,
		0x0,
		0x20202020200,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x402010080400,
		0x0,
		0x2020202020200,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x2),
		0x0,
		0x0,
		0x0,
		0x8,
		0x18,
		0x38,
		0x78,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x200,
		0x0,
		0x400,
		0x0,
		0x800,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40400,
		0x0,
		0x0,
		0x100800,
		0x0,
		0x0,
		0x0,
		0x0,
		0x4040400,
		0x0,
		0x0,
		0x0,
		0x20100800,
		0x0,
		0x0,
		0x0,
		0x404040400,
		0x0,
		0x0,
		0x0,
		0x0,
		0x4020100800,
		0x0,
		0x0,
		0x40404040400,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x4040404040400,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x6),
		0x4,
		0x0,
		0x0,
		0x0,
		0x10,
		0x30,
		0x70,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x400,
		0x0,
		0x800,
		0x0,
		0x1000,
		0x0,
		0x0,
		0x20400,
		0x0,
		0x0,
		0x80800,
		0x0,
		0x0,
		0x201000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x8080800,
		0x0,
		0x0,
		0x0,
		0x40201000,
		0x0,
		0x0,
		0x0,
		0x808080800,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x80808080800,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x8080808080800,
		0x0,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0xE),
		0xC,
		0x8,
		0x0,
		0x0,
		0x0,
		0x20,
		0x60,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x800,
		0x0,
		0x1000,
		0x0,
		0x2000,
		0x0,
		0x0,
		0x40800,
		0x0,
		0x0,
		0x101000,
		0x0,
		0x0,
		0x402000,
		0x2040800,
		0x0,
		0x0,
		0x0,
		0x10101000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x1010101000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x101010101000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x10101010101000,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x1E),
		0x1C,
		0x18,
		0x10,
		0x0,
		0x0,
		0x0,
		0x40,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x1000,
		0x0,
		0x2000,
		0x0,
		0x4000,
		0x0,
		0x0,
		0x81000,
		0x0,
		0x0,
		0x202000,
		0x0,
		0x0,
		0x0,
		0x4081000,
		0x0,
		0x0,
		0x0,
		0x20202000,
		0x0,
		0x0,
		0x204081000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2020202000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x202020202000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20202020202000,
		0x0,
		0x0,
	],
	[
		Bitboard(0x3E),
		0x3C,
		0x38,
		0x30,
		0x20,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2000,
		0x0,
		0x4000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x102000,
		0x0,
		0x0,
		0x404000,
		0x0,
		0x0,
		0x0,
		0x8102000,
		0x0,
		0x0,
		0x0,
		0x40404000,
		0x0,
		0x0,
		0x408102000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x4040404000,
		0x0,
		0x20408102000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x404040404000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40404040404000,
		0x0,
	],
	[
		Bitboard(0x7E),
		0x7C,
		0x78,
		0x70,
		0x60,
		0x40,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x4000,
		0x0,
		0x8000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x204000,
		0x0,
		0x0,
		0x808000,
		0x0,
		0x0,
		0x0,
		0x10204000,
		0x0,
		0x0,
		0x0,
		0x80808000,
		0x0,
		0x0,
		0x810204000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x8080808000,
		0x0,
		0x40810204000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x808080808000,
		0x2040810204000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x80808080808000,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x200,
		0x600,
		0xE00,
		0x1E00,
		0x3E00,
		0x7E00,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x10000,
		0x0,
		0x20000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x1010000,
		0x0,
		0x0,
		0x4020000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x101010000,
		0x0,
		0x0,
		0x0,
		0x804020000,
		0x0,
		0x0,
		0x0,
		0x10101010000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x100804020000,
		0x0,
		0x0,
		0x1010101010000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20100804020000,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x400,
		0xC00,
		0x1C00,
		0x3C00,
		0x7C00,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20000,
		0x0,
		0x40000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2020000,
		0x0,
		0x0,
		0x8040000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x202020000,
		0x0,
		0x0,
		0x0,
		0x1008040000,
		0x0,
		0x0,
		0x0,
		0x20202020000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x201008040000,
		0x0,
		0x0,
		0x2020202020000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40201008040000,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x200,
		0x0,
		0x0,
		0x0,
		0x800,
		0x1800,
		0x3800,
		0x7800,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20000,
		0x0,
		0x40000,
		0x0,
		0x80000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x4040000,
		0x0,
		0x0,
		0x10080000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x404040000,
		0x0,
		0x0,
		0x0,
		0x2010080000,
		0x0,
		0x0,
		0x0,
		0x40404040000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x402010080000,
		0x0,
		0x0,
		0x4040404040000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x600,
		0x400,
		0x0,
		0x0,
		0x0,
		0x1000,
		0x3000,
		0x7000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40000,
		0x0,
		0x80000,
		0x0,
		0x100000,
		0x0,
		0x0,
		0x2040000,
		0x0,
		0x0,
		0x8080000,
		0x0,
		0x0,
		0x20100000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x808080000,
		0x0,
		0x0,
		0x0,
		0x4020100000,
		0x0,
		0x0,
		0x0,
		0x80808080000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x8080808080000,
		0x0,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0xE00,
		0xC00,
		0x800,
		0x0,
		0x0,
		0x0,
		0x2000,
		0x6000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x80000,
		0x0,
		0x100000,
		0x0,
		0x200000,
		0x0,
		0x0,
		0x4080000,
		0x0,
		0x0,
		0x10100000,
		0x0,
		0x0,
		0x40200000,
		0x204080000,
		0x0,
		0x0,
		0x0,
		0x1010100000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x101010100000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x10101010100000,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x1E00,
		0x1C00,
		0x1800,
		0x1000,
		0x0,
		0x0,
		0x0,
		0x4000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x100000,
		0x0,
		0x200000,
		0x0,
		0x400000,
		0x0,
		0x0,
		0x8100000,
		0x0,
		0x0,
		0x20200000,
		0x0,
		0x0,
		0x0,
		0x408100000,
		0x0,
		0x0,
		0x0,
		0x2020200000,
		0x0,
		0x0,
		0x20408100000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x202020200000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20202020200000,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x3E00,
		0x3C00,
		0x3800,
		0x3000,
		0x2000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x200000,
		0x0,
		0x400000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x10200000,
		0x0,
		0x0,
		0x40400000,
		0x0,
		0x0,
		0x0,
		0x810200000,
		0x0,
		0x0,
		0x0,
		0x4040400000,
		0x0,
		0x0,
		0x40810200000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x404040400000,
		0x0,
		0x2040810200000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40404040400000,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x7E00,
		0x7C00,
		0x7800,
		0x7000,
		0x6000,
		0x4000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x400000,
		0x0,
		0x800000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20400000,
		0x0,
		0x0,
		0x80800000,
		0x0,
		0x0,
		0x0,
		0x1020400000,
		0x0,
		0x0,
		0x0,
		0x8080800000,
		0x0,
		0x0,
		0x81020400000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x808080800000,
		0x0,
		0x4081020400000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x80808080800000,
	],
	[
		Bitboard(0x100),
		0x0,
		0x200,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20000,
		0x60000,
		0xE0000,
		0x1E0000,
		0x3E0000,
		0x7E0000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x1000000,
		0x0,
		0x2000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x101000000,
		0x0,
		0x0,
		0x402000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x10101000000,
		0x0,
		0x0,
		0x0,
		0x80402000000,
		0x0,
		0x0,
		0x0,
		0x1010101000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x10080402000000,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x200,
		0x0,
		0x400,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40000,
		0xC0000,
		0x1C0000,
		0x3C0000,
		0x7C0000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2000000,
		0x0,
		0x4000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x202000000,
		0x0,
		0x0,
		0x804000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20202000000,
		0x0,
		0x0,
		0x0,
		0x100804000000,
		0x0,
		0x0,
		0x0,
		0x2020202000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20100804000000,
		0x0,
	],
	[
		Bitboard(0x200),
		0x0,
		0x400,
		0x0,
		0x800,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20000,
		0x0,
		0x0,
		0x0,
		0x80000,
		0x180000,
		0x380000,
		0x780000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2000000,
		0x0,
		0x4000000,
		0x0,
		0x8000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x404000000,
		0x0,
		0x0,
		0x1008000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40404000000,
		0x0,
		0x0,
		0x0,
		0x201008000000,
		0x0,
		0x0,
		0x0,
		0x4040404000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40201008000000,
	],
	[
		Bitboard(0x0),
		0x400,
		0x0,
		0x800,
		0x0,
		0x1000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x60000,
		0x40000,
		0x0,
		0x0,
		0x0,
		0x100000,
		0x300000,
		0x700000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x4000000,
		0x0,
		0x8000000,
		0x0,
		0x10000000,
		0x0,
		0x0,
		0x204000000,
		0x0,
		0x0,
		0x808000000,
		0x0,
		0x0,
		0x2010000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x80808000000,
		0x0,
		0x0,
		0x0,
		0x402010000000,
		0x0,
		0x0,
		0x0,
		0x8080808000000,
		0x0,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x800,
		0x0,
		0x1000,
		0x0,
		0x2000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0xE0000,
		0xC0000,
		0x80000,
		0x0,
		0x0,
		0x0,
		0x200000,
		0x600000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x8000000,
		0x0,
		0x10000000,
		0x0,
		0x20000000,
		0x0,
		0x0,
		0x408000000,
		0x0,
		0x0,
		0x1010000000,
		0x0,
		0x0,
		0x4020000000,
		0x20408000000,
		0x0,
		0x0,
		0x0,
		0x101010000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x10101010000000,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x1000,
		0x0,
		0x2000,
		0x0,
		0x4000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x1E0000,
		0x1C0000,
		0x180000,
		0x100000,
		0x0,
		0x0,
		0x0,
		0x400000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x10000000,
		0x0,
		0x20000000,
		0x0,
		0x40000000,
		0x0,
		0x0,
		0x810000000,
		0x0,
		0x0,
		0x2020000000,
		0x0,
		0x0,
		0x0,
		0x40810000000,
		0x0,
		0x0,
		0x0,
		0x202020000000,
		0x0,
		0x0,
		0x2040810000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20202020000000,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x0,
		0x2000,
		0x0,
		0x4000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x3E0000,
		0x3C0000,
		0x380000,
		0x300000,
		0x200000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20000000,
		0x0,
		0x40000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x1020000000,
		0x0,
		0x0,
		0x4040000000,
		0x0,
		0x0,
		0x0,
		0x81020000000,
		0x0,
		0x0,
		0x0,
		0x404040000000,
		0x0,
		0x0,
		0x4081020000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40404040000000,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x0,
		0x0,
		0x4000,
		0x0,
		0x8000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x7E0000,
		0x7C0000,
		0x780000,
		0x700000,
		0x600000,
		0x400000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40000000,
		0x0,
		0x80000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2040000000,
		0x0,
		0x0,
		0x8080000000,
		0x0,
		0x0,
		0x0,
		0x102040000000,
		0x0,
		0x0,
		0x0,
		0x808080000000,
		0x0,
		0x0,
		0x8102040000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x80808080000000,
	],
	[
		Bitboard(0x10100),
		0x0,
		0x0,
		0x20400,
		0x0,
		0x0,
		0x0,
		0x0,
		0x10000,
		0x0,
		0x20000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2000000,
		0x6000000,
		0xE000000,
		0x1E000000,
		0x3E000000,
		0x7E000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x100000000,
		0x0,
		0x200000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x10100000000,
		0x0,
		0x0,
		0x40200000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x1010100000000,
		0x0,
		0x0,
		0x0,
		0x8040200000000,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x20200,
		0x0,
		0x0,
		0x40800,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20000,
		0x0,
		0x40000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x4000000,
		0xC000000,
		0x1C000000,
		0x3C000000,
		0x7C000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x200000000,
		0x0,
		0x400000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20200000000,
		0x0,
		0x0,
		0x80400000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2020200000000,
		0x0,
		0x0,
		0x0,
		0x10080400000000,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x40400,
		0x0,
		0x0,
		0x81000,
		0x0,
		0x0,
		0x20000,
		0x0,
		0x40000,
		0x0,
		0x80000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2000000,
		0x0,
		0x0,
		0x0,
		0x8000000,
		0x18000000,
		0x38000000,
		0x78000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x200000000,
		0x0,
		0x400000000,
		0x0,
		0x800000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40400000000,
		0x0,
		0x0,
		0x100800000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x4040400000000,
		0x0,
		0x0,
		0x0,
		0x20100800000000,
		0x0,
	],
	[
		Bitboard(0x40200),
		0x0,
		0x0,
		0x80800,
		0x0,
		0x0,
		0x102000,
		0x0,
		0x0,
		0x40000,
		0x0,
		0x80000,
		0x0,
		0x100000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x6000000,
		0x4000000,
		0x0,
		0x0,
		0x0,
		0x10000000,
		0x30000000,
		0x70000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x400000000,
		0x0,
		0x800000000,
		0x0,
		0x1000000000,
		0x0,
		0x0,
		0x20400000000,
		0x0,
		0x0,
		0x80800000000,
		0x0,
		0x0,
		0x201000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x8080800000000,
		0x0,
		0x0,
		0x0,
		0x40201000000000,
	],
	[
		Bitboard(0x0),
		0x80400,
		0x0,
		0x0,
		0x101000,
		0x0,
		0x0,
		0x204000,
		0x0,
		0x0,
		0x80000,
		0x0,
		0x100000,
		0x0,
		0x200000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0xE000000,
		0xC000000,
		0x8000000,
		0x0,
		0x0,
		0x0,
		0x20000000,
		0x60000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x800000000,
		0x0,
		0x1000000000,
		0x0,
		0x2000000000,
		0x0,
		0x0,
		0x40800000000,
		0x0,
		0x0,
		0x101000000000,
		0x0,
		0x0,
		0x402000000000,
		0x2040800000000,
		0x0,
		0x0,
		0x0,
		0x10101000000000,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x100800,
		0x0,
		0x0,
		0x202000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x100000,
		0x0,
		0x200000,
		0x0,
		0x400000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x1E000000,
		0x1C000000,
		0x18000000,
		0x10000000,
		0x0,
		0x0,
		0x0,
		0x40000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x1000000000,
		0x0,
		0x2000000000,
		0x0,
		0x4000000000,
		0x0,
		0x0,
		0x81000000000,
		0x0,
		0x0,
		0x202000000000,
		0x0,
		0x0,
		0x0,
		0x4081000000000,
		0x0,
		0x0,
		0x0,
		0x20202000000000,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x201000,
		0x0,
		0x0,
		0x404000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x200000,
		0x0,
		0x400000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x3E000000,
		0x3C000000,
		0x38000000,
		0x30000000,
		0x20000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2000000000,
		0x0,
		0x4000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x102000000000,
		0x0,
		0x0,
		0x404000000000,
		0x0,
		0x0,
		0x0,
		0x8102000000000,
		0x0,
		0x0,
		0x0,
		0x40404000000000,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x0,
		0x402000,
		0x0,
		0x0,
		0x808000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x400000,
		0x0,
		0x800000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x7E000000,
		0x7C000000,
		0x78000000,
		0x70000000,
		0x60000000,
		0x40000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x4000000000,
		0x0,
		0x8000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x204000000000,
		0x0,
		0x0,
		0x808000000000,
		0x0,
		0x0,
		0x0,
		0x10204000000000,
		0x0,
		0x0,
		0x0,
		0x80808000000000,
	],
	[
		Bitboard(0x1010100),
		0x0,
		0x0,
		0x0,
		0x2040800,
		0x0,
		0x0,
		0x0,
		0x1010000,
		0x0,
		0x0,
		0x2040000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x1000000,
		0x0,
		0x2000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x200000000,
		0x600000000,
		0xE00000000,
		0x1E00000000,
		0x3E00000000,
		0x7E00000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x10000000000,
		0x0,
		0x20000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x1010000000000,
		0x0,
		0x0,
		0x4020000000000,
		0x0,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x2020200,
		0x0,
		0x0,
		0x0,
		0x4081000,
		0x0,
		0x0,
		0x0,
		0x2020000,
		0x0,
		0x0,
		0x4080000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2000000,
		0x0,
		0x4000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x400000000,
		0xC00000000,
		0x1C00000000,
		0x3C00000000,
		0x7C00000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20000000000,
		0x0,
		0x40000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2020000000000,
		0x0,
		0x0,
		0x8040000000000,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x4040400,
		0x0,
		0x0,
		0x0,
		0x8102000,
		0x0,
		0x0,
		0x0,
		0x4040000,
		0x0,
		0x0,
		0x8100000,
		0x0,
		0x0,
		0x2000000,
		0x0,
		0x4000000,
		0x0,
		0x8000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x200000000,
		0x0,
		0x0,
		0x0,
		0x800000000,
		0x1800000000,
		0x3800000000,
		0x7800000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20000000000,
		0x0,
		0x40000000000,
		0x0,
		0x80000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x4040000000000,
		0x0,
		0x0,
		0x10080000000000,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x8080800,
		0x0,
		0x0,
		0x0,
		0x10204000,
		0x4020000,
		0x0,
		0x0,
		0x8080000,
		0x0,
		0x0,
		0x10200000,
		0x0,
		0x0,
		0x4000000,
		0x0,
		0x8000000,
		0x0,
		0x10000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x600000000,
		0x400000000,
		0x0,
		0x0,
		0x0,
		0x1000000000,
		0x3000000000,
		0x7000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40000000000,
		0x0,
		0x80000000000,
		0x0,
		0x100000000000,
		0x0,
		0x0,
		0x2040000000000,
		0x0,
		0x0,
		0x8080000000000,
		0x0,
		0x0,
		0x20100000000000,
		0x0,
	],
	[
		Bitboard(0x8040200),
		0x0,
		0x0,
		0x0,
		0x10101000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x8040000,
		0x0,
		0x0,
		0x10100000,
		0x0,
		0x0,
		0x20400000,
		0x0,
		0x0,
		0x8000000,
		0x0,
		0x10000000,
		0x0,
		0x20000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0xE00000000,
		0xC00000000,
		0x800000000,
		0x0,
		0x0,
		0x0,
		0x2000000000,
		0x6000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x80000000000,
		0x0,
		0x100000000000,
		0x0,
		0x200000000000,
		0x0,
		0x0,
		0x4080000000000,
		0x0,
		0x0,
		0x10100000000000,
		0x0,
		0x0,
		0x40200000000000,
	],
	[
		Bitboard(0x0),
		0x10080400,
		0x0,
		0x0,
		0x0,
		0x20202000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x10080000,
		0x0,
		0x0,
		0x20200000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x10000000,
		0x0,
		0x20000000,
		0x0,
		0x40000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x1E00000000,
		0x1C00000000,
		0x1800000000,
		0x1000000000,
		0x0,
		0x0,
		0x0,
		0x4000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x100000000000,
		0x0,
		0x200000000000,
		0x0,
		0x400000000000,
		0x0,
		0x0,
		0x8100000000000,
		0x0,
		0x0,
		0x20200000000000,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x20100800,
		0x0,
		0x0,
		0x0,
		0x40404000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20100000,
		0x0,
		0x0,
		0x40400000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20000000,
		0x0,
		0x40000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x3E00000000,
		0x3C00000000,
		0x3800000000,
		0x3000000000,
		0x2000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x200000000000,
		0x0,
		0x400000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x10200000000000,
		0x0,
		0x0,
		0x40400000000000,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x40201000,
		0x0,
		0x0,
		0x0,
		0x80808000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40200000,
		0x0,
		0x0,
		0x80800000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40000000,
		0x0,
		0x80000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x7E00000000,
		0x7C00000000,
		0x7800000000,
		0x7000000000,
		0x6000000000,
		0x4000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x400000000000,
		0x0,
		0x800000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20400000000000,
		0x0,
		0x0,
		0x80800000000000,
	],
	[
		Bitboard(0x101010100),
		0x0,
		0x0,
		0x0,
		0x0,
		0x204081000,
		0x0,
		0x0,
		0x101010000,
		0x0,
		0x0,
		0x0,
		0x204080000,
		0x0,
		0x0,
		0x0,
		0x101000000,
		0x0,
		0x0,
		0x204000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x100000000,
		0x0,
		0x200000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20000000000,
		0x60000000000,
		0xE0000000000,
		0x1E0000000000,
		0x3E0000000000,
		0x7E0000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x1000000000000,
		0x0,
		0x2000000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x202020200,
		0x0,
		0x0,
		0x0,
		0x0,
		0x408102000,
		0x0,
		0x0,
		0x202020000,
		0x0,
		0x0,
		0x0,
		0x408100000,
		0x0,
		0x0,
		0x0,
		0x202000000,
		0x0,
		0x0,
		0x408000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x200000000,
		0x0,
		0x400000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40000000000,
		0xC0000000000,
		0x1C0000000000,
		0x3C0000000000,
		0x7C0000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2000000000000,
		0x0,
		0x4000000000000,
		0x0,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x404040400,
		0x0,
		0x0,
		0x0,
		0x0,
		0x810204000,
		0x0,
		0x0,
		0x404040000,
		0x0,
		0x0,
		0x0,
		0x810200000,
		0x0,
		0x0,
		0x0,
		0x404000000,
		0x0,
		0x0,
		0x810000000,
		0x0,
		0x0,
		0x200000000,
		0x0,
		0x400000000,
		0x0,
		0x800000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20000000000,
		0x0,
		0x0,
		0x0,
		0x80000000000,
		0x180000000000,
		0x380000000000,
		0x780000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2000000000000,
		0x0,
		0x4000000000000,
		0x0,
		0x8000000000000,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x808080800,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x808080000,
		0x0,
		0x0,
		0x0,
		0x1020400000,
		0x402000000,
		0x0,
		0x0,
		0x808000000,
		0x0,
		0x0,
		0x1020000000,
		0x0,
		0x0,
		0x400000000,
		0x0,
		0x800000000,
		0x0,
		0x1000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x60000000000,
		0x40000000000,
		0x0,
		0x0,
		0x0,
		0x100000000000,
		0x300000000000,
		0x700000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x4000000000000,
		0x0,
		0x8000000000000,
		0x0,
		0x10000000000000,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x0,
		0x1010101000,
		0x0,
		0x0,
		0x0,
		0x804020000,
		0x0,
		0x0,
		0x0,
		0x1010100000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x804000000,
		0x0,
		0x0,
		0x1010000000,
		0x0,
		0x0,
		0x2040000000,
		0x0,
		0x0,
		0x800000000,
		0x0,
		0x1000000000,
		0x0,
		0x2000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0xE0000000000,
		0xC0000000000,
		0x80000000000,
		0x0,
		0x0,
		0x0,
		0x200000000000,
		0x600000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x8000000000000,
		0x0,
		0x10000000000000,
		0x0,
		0x20000000000000,
		0x0,
	],
	[
		Bitboard(0x1008040200),
		0x0,
		0x0,
		0x0,
		0x0,
		0x2020202000,
		0x0,
		0x0,
		0x0,
		0x1008040000,
		0x0,
		0x0,
		0x0,
		0x2020200000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x1008000000,
		0x0,
		0x0,
		0x2020000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x1000000000,
		0x0,
		0x2000000000,
		0x0,
		0x4000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x1E0000000000,
		0x1C0000000000,
		0x180000000000,
		0x100000000000,
		0x0,
		0x0,
		0x0,
		0x400000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x10000000000000,
		0x0,
		0x20000000000000,
		0x0,
		0x40000000000000,
	],
	[
		Bitboard(0x0),
		0x2010080400,
		0x0,
		0x0,
		0x0,
		0x0,
		0x4040404000,
		0x0,
		0x0,
		0x0,
		0x2010080000,
		0x0,
		0x0,
		0x0,
		0x4040400000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2010000000,
		0x0,
		0x0,
		0x4040000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2000000000,
		0x0,
		0x4000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x3E0000000000,
		0x3C0000000000,
		0x380000000000,
		0x300000000000,
		0x200000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20000000000000,
		0x0,
		0x40000000000000,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x4020100800,
		0x0,
		0x0,
		0x0,
		0x0,
		0x8080808000,
		0x0,
		0x0,
		0x0,
		0x4020100000,
		0x0,
		0x0,
		0x0,
		0x8080800000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x4020000000,
		0x0,
		0x0,
		0x8080000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x4000000000,
		0x0,
		0x8000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x7E0000000000,
		0x7C0000000000,
		0x780000000000,
		0x700000000000,
		0x600000000000,
		0x400000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40000000000000,
		0x0,
		0x80000000000000,
	],
	[
		Bitboard(0x10101010100),
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20408102000,
		0x0,
		0x10101010000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20408100000,
		0x0,
		0x0,
		0x10101000000,
		0x0,
		0x0,
		0x0,
		0x20408000000,
		0x0,
		0x0,
		0x0,
		0x10100000000,
		0x0,
		0x0,
		0x20400000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x10000000000,
		0x0,
		0x20000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2000000000000,
		0x6000000000000,
		0xE000000000000,
		0x1E000000000000,
		0x3E000000000000,
		0x7E000000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x20202020200,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40810204000,
		0x0,
		0x20202020000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40810200000,
		0x0,
		0x0,
		0x20202000000,
		0x0,
		0x0,
		0x0,
		0x40810000000,
		0x0,
		0x0,
		0x0,
		0x20200000000,
		0x0,
		0x0,
		0x40800000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20000000000,
		0x0,
		0x40000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x4000000000000,
		0xC000000000000,
		0x1C000000000000,
		0x3C000000000000,
		0x7C000000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x40404040400,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40404040000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x81020400000,
		0x0,
		0x0,
		0x40404000000,
		0x0,
		0x0,
		0x0,
		0x81020000000,
		0x0,
		0x0,
		0x0,
		0x40400000000,
		0x0,
		0x0,
		0x81000000000,
		0x0,
		0x0,
		0x20000000000,
		0x0,
		0x40000000000,
		0x0,
		0x80000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2000000000000,
		0x0,
		0x0,
		0x0,
		0x8000000000000,
		0x18000000000000,
		0x38000000000000,
		0x78000000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x80808080800,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x80808080000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x80808000000,
		0x0,
		0x0,
		0x0,
		0x102040000000,
		0x40200000000,
		0x0,
		0x0,
		0x80800000000,
		0x0,
		0x0,
		0x102000000000,
		0x0,
		0x0,
		0x40000000000,
		0x0,
		0x80000000000,
		0x0,
		0x100000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x6000000000000,
		0x4000000000000,
		0x0,
		0x0,
		0x0,
		0x10000000000000,
		0x30000000000000,
		0x70000000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x0,
		0x101010101000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x101010100000,
		0x0,
		0x0,
		0x0,
		0x80402000000,
		0x0,
		0x0,
		0x0,
		0x101010000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x80400000000,
		0x0,
		0x0,
		0x101000000000,
		0x0,
		0x0,
		0x204000000000,
		0x0,
		0x0,
		0x80000000000,
		0x0,
		0x100000000000,
		0x0,
		0x200000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0xE000000000000,
		0xC000000000000,
		0x8000000000000,
		0x0,
		0x0,
		0x0,
		0x20000000000000,
		0x60000000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x0,
		0x0,
		0x202020202000,
		0x0,
		0x0,
		0x100804020000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x202020200000,
		0x0,
		0x0,
		0x0,
		0x100804000000,
		0x0,
		0x0,
		0x0,
		0x202020000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x100800000000,
		0x0,
		0x0,
		0x202000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x100000000000,
		0x0,
		0x200000000000,
		0x0,
		0x400000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x1E000000000000,
		0x1C000000000000,
		0x18000000000000,
		0x10000000000000,
		0x0,
		0x0,
		0x0,
		0x40000000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x201008040200),
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x404040404000,
		0x0,
		0x0,
		0x201008040000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x404040400000,
		0x0,
		0x0,
		0x0,
		0x201008000000,
		0x0,
		0x0,
		0x0,
		0x404040000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x201000000000,
		0x0,
		0x0,
		0x404000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x200000000000,
		0x0,
		0x400000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x3E000000000000,
		0x3C000000000000,
		0x38000000000000,
		0x30000000000000,
		0x20000000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x0),
		0x402010080400,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x808080808000,
		0x0,
		0x0,
		0x402010080000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x808080800000,
		0x0,
		0x0,
		0x0,
		0x402010000000,
		0x0,
		0x0,
		0x0,
		0x808080000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x402000000000,
		0x0,
		0x0,
		0x808000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x400000000000,
		0x0,
		0x800000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x7E000000000000,
		0x7C000000000000,
		0x78000000000000,
		0x70000000000000,
		0x60000000000000,
		0x40000000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x1010101010100),
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2040810204000,
		0x1010101010000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2040810200000,
		0x0,
		0x1010101000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2040810000000,
		0x0,
		0x0,
		0x1010100000000,
		0x0,
		0x0,
		0x0,
		0x2040800000000,
		0x0,
		0x0,
		0x0,
		0x1010000000000,
		0x0,
		0x0,
		0x2040000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x1000000000000,
		0x0,
		0x2000000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x200000000000000,
		0x600000000000000,
		0xE00000000000000,
		0x1E00000000000000,
		0x3E00000000000000,
		0x7E00000000000000,
	],
	[
		Bitboard(0x0),
		0x2020202020200,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2020202020000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x4081020400000,
		0x0,
		0x2020202000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x4081020000000,
		0x0,
		0x0,
		0x2020200000000,
		0x0,
		0x0,
		0x0,
		0x4081000000000,
		0x0,
		0x0,
		0x0,
		0x2020000000000,
		0x0,
		0x0,
		0x4080000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x2000000000000,
		0x0,
		0x4000000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x400000000000000,
		0xC00000000000000,
		0x1C00000000000000,
		0x3C00000000000000,
		0x7C00000000000000,
	],
	[
		Bitboard(0x0),
		0x0,
		0x4040404040400,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x4040404040000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x4040404000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x8102040000000,
		0x0,
		0x0,
		0x4040400000000,
		0x0,
		0x0,
		0x0,
		0x8102000000000,
		0x0,
		0x0,
		0x0,
		0x4040000000000,
		0x0,
		0x0,
		0x8100000000000,
		0x0,
		0x0,
		0x2000000000000,
		0x0,
		0x4000000000000,
		0x0,
		0x8000000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x200000000000000,
		0x0,
		0x0,
		0x0,
		0x800000000000000,
		0x1800000000000000,
		0x3800000000000000,
		0x7800000000000000,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x8080808080800,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x8080808080000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x8080808000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x8080800000000,
		0x0,
		0x0,
		0x0,
		0x10204000000000,
		0x4020000000000,
		0x0,
		0x0,
		0x8080000000000,
		0x0,
		0x0,
		0x10200000000000,
		0x0,
		0x0,
		0x4000000000000,
		0x0,
		0x8000000000000,
		0x0,
		0x10000000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x600000000000000,
		0x400000000000000,
		0x0,
		0x0,
		0x0,
		0x1000000000000000,
		0x3000000000000000,
		0x7000000000000000,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x0,
		0x10101010101000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x10101010100000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x10101010000000,
		0x0,
		0x0,
		0x0,
		0x8040200000000,
		0x0,
		0x0,
		0x0,
		0x10101000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x8040000000000,
		0x0,
		0x0,
		0x10100000000000,
		0x0,
		0x0,
		0x20400000000000,
		0x0,
		0x0,
		0x8000000000000,
		0x0,
		0x10000000000000,
		0x0,
		0x20000000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0xE00000000000000,
		0xC00000000000000,
		0x800000000000000,
		0x0,
		0x0,
		0x0,
		0x2000000000000000,
		0x6000000000000000,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x0,
		0x0,
		0x20202020202000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20202020200000,
		0x0,
		0x0,
		0x10080402000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20202020000000,
		0x0,
		0x0,
		0x0,
		0x10080400000000,
		0x0,
		0x0,
		0x0,
		0x20202000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x10080000000000,
		0x0,
		0x0,
		0x20200000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x10000000000000,
		0x0,
		0x20000000000000,
		0x0,
		0x40000000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x1E00000000000000,
		0x1C00000000000000,
		0x1800000000000000,
		0x1000000000000000,
		0x0,
		0x0,
		0x0,
		0x4000000000000000,
	],
	[
		Bitboard(0x0),
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40404040404000,
		0x0,
		0x20100804020000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40404040400000,
		0x0,
		0x0,
		0x20100804000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40404040000000,
		0x0,
		0x0,
		0x0,
		0x20100800000000,
		0x0,
		0x0,
		0x0,
		0x40404000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20100000000000,
		0x0,
		0x0,
		0x40400000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x20000000000000,
		0x0,
		0x40000000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x3E00000000000000,
		0x3C00000000000000,
		0x3800000000000000,
		0x3000000000000000,
		0x2000000000000000,
		0x0,
		0x0,
		0x0,
	],
	[
		Bitboard(0x40201008040200),
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x80808080808000,
		0x0,
		0x40201008040000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x80808080800000,
		0x0,
		0x0,
		0x40201008000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x80808080000000,
		0x0,
		0x0,
		0x0,
		0x40201000000000,
		0x0,
		0x0,
		0x0,
		0x80808000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40200000000000,
		0x0,
		0x0,
		0x80800000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x40000000000000,
		0x0,
		0x80000000000000,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x0,
		0x7E00000000000000,
		0x7C00000000000000,
		0x7800000000000000,
		0x7000000000000000,
		0x6000000000000000,
		0x4000000000000000,
		0x0,
		0x0,
	],
]