module engine

pub struct EngineInfo {
pub:
	name    string = 'Visionary IX'
	version string = '0.2.1'
	author  string = 'tabledotnet'
}
