module engine

pub struct EngineInfo {
pub:
	name    string = 'Visionary IX'
	version string = '0.5'
	author  string = 'tabledotnet'
}
