module chess

pub const bishop_magics = [
        Magic { 0x40201008040200, 0x1004600204002280, 58, 0 },
        Magic { 0x402010080400, 0x20220400608004, 59, 64 },
        Magic { 0x4020100A00, 0x4440092041001, 59, 96 },
        Magic { 0x40221400, 0x6048204840109080, 59, 128 },
        Magic { 0x2442800, 0x2021010108943, 59, 160 },
        Magic { 0x204085000, 0xA400822020080030, 59, 192 },
        Magic { 0x20408102000, 0x80C808888400400, 59, 224 },
        Magic { 0x2040810204000, 0x8000220800880900, 58, 256 },
        Magic { 0x20100804020000, 0x4A80180810040842, 59, 320 },
        Magic { 0x40201008040000, 0x30240404044200, 59, 352 },
        Magic { 0x4020100A0000, 0x424202002002, 59, 384 },
        Magic { 0x4022140000, 0x1000109082080008, 59, 416 },
        Magic { 0x244280000, 0x802508820400000, 59, 448 },
        Magic { 0x20408500000, 0x103A920802180444, 59, 480 },
        Magic { 0x2040810200000, 0x4000008188084022, 59, 512 },
        Magic { 0x4081020400000, 0xB000C1C8080802, 59, 544 },
        Magic { 0x10080402000200, 0x4140040808810402, 59, 576 },
        Magic { 0x20100804000400, 0x308010210A40580, 59, 608 },
        Magic { 0x4020100A000A00, 0x900001810E0020, 57, 640 },
        Magic { 0x402214001400, 0x8008402142040, 57, 768 },
        Magic { 0x24428002800, 0x141000820080010, 57, 896 },
        Magic { 0x2040850005000, 0x4006010822032000, 57, 1024 },
        Magic { 0x4081020002000, 0x400809048183801, 59, 1152 },
        Magic { 0x8102040004000, 0x905001044020141, 59, 1184 },
        Magic { 0x8040200020400, 0x20040008703400, 59, 1216 },
        Magic { 0x10080400040800, 0x1108240002040800, 59, 1248 },
        Magic { 0x20100A000A1000, 0x1044240062040408, 57, 1280 },
        Magic { 0x40221400142200, 0x2840401C010200, 55, 1408 },
        Magic { 0x2442800284400, 0x2848800C002000, 55, 1920 },
        Magic { 0x4085000500800, 0x8004010008104202, 57, 2432 },
        Magic { 0x8102000201000, 0xD011200044A1000, 59, 2560 },
        Magic { 0x10204000402000, 0x4004000806410, 59, 2592 },
        Magic { 0x4020002040800, 0x24042458202100, 59, 2624 },
        Magic { 0x8040004081000, 0x2188040210100200, 59, 2656 },
        Magic { 0x100A000A102000, 0x808404044081A0, 57, 2688 },
        Magic { 0x22140014224000, 0x651020081180080, 55, 2816 },
        Magic { 0x44280028440200, 0x40420400C20108, 55, 3328 },
        Magic { 0x8500050080400, 0x384040090080802, 57, 3840 },
        Magic { 0x10200020100800, 0x148A80280064200, 59, 3968 },
        Magic { 0x20400040201000, 0x1814011A0010C241, 59, 4000 },
        Magic { 0x2000204081000, 0x8008021050081410, 59, 4032 },
        Magic { 0x4000408102000, 0xA080128415410, 59, 4064 },
        Magic { 0xA000A10204000, 0x220280280800C100, 57, 4096 },
        Magic { 0x14001422400000, 0x40002018000102, 57, 4224 },
        Magic { 0x28002844020000, 0x400100200640200, 57, 4352 },
        Magic { 0x50005008040200, 0x21102302004140, 57, 4480 },
        Magic { 0x20002010080400, 0x60012212020080, 59, 4608 },
        Magic { 0x40004020100800, 0x200442808104420E, 59, 4640 },
        Magic { 0x20408102000, 0x144453010100800, 59, 4672 },
        Magic { 0x40810204000, 0x21050110520200, 59, 4704 },
        Magic { 0xA1020400000, 0x100804442C040040, 59, 4736 },
        Magic { 0x142240000000, 0x4000002020882200, 59, 4768 },
        Magic { 0x284402000000, 0x100200400A820141, 59, 4800 },
        Magic { 0x500804020000, 0x1A00400801010410, 59, 4832 },
        Magic { 0x201008040200, 0x10208802808010, 59, 4864 },
        Magic { 0x402010080400, 0x20080100408021, 59, 4896 },
        Magic { 0x2040810204000, 0x2010048040400, 58, 4928 },
        Magic { 0x4081020400000, 0x9008214402080301, 59, 4992 },
        Magic { 0xA102040000000, 0x40300062A011020, 59, 5024 },
        Magic { 0x14224000000000, 0x38130801420204, 59, 5056 },
        Magic { 0x28440200000000, 0x2402A8034504C00, 59, 5088 },
        Magic { 0x50080402000000, 0x900012014410201, 59, 5120 },
        Magic { 0x20100804020000, 0x1410A0C012200, 59, 5152 },
        Magic { 0x40201008040200, 0x4011013904040040, 58, 5184 },
]
pub const bishop_table_size = 5248

pub const rook_magics = [
        Magic { 0x101010101017E, 0x80002040028018, 52, 0 },
        Magic { 0x202020202027E, 0x4081040200110, 52, 4096 },
        Magic { 0x404040404047E, 0x2500080460001040, 52, 8192 },
        Magic { 0x808080808087E, 0x780040210002800, 52, 12288 },
        Magic { 0x1010101010107E, 0x280040008000182, 52, 16384 },
        Magic { 0x2020202020207E, 0x2B00020804004081, 52, 20480 },
        Magic { 0x4040404040407E, 0x400004094100802, 52, 24576 },
        Magic { 0x8080808080807E, 0x480002040800100, 52, 28672 },
        Magic { 0x1010101017F00, 0x5012800022400210, 52, 32768 },
        Magic { 0x2020202027C00, 0x2122804000892000, 54, 36864 },
        Magic { 0x4040404047A00, 0x801000806003, 54, 37888 },
        Magic { 0x8080808087600, 0xC128801000800801, 54, 38912 },
        Magic { 0x10101010106E00, 0x28070011005800C4, 54, 39936 },
        Magic { 0x20202020205E00, 0x48A000408820010, 54, 40960 },
        Magic { 0x40404040403E00, 0x9200AA00050804, 54, 41984 },
        Magic { 0x8080808080FE00, 0x9000180A20151, 52, 43008 },
        Magic { 0x10101017F0100, 0x2828D08000400028, 52, 47104 },
        Magic { 0x20202027C0200, 0x1150A0022008042, 54, 51200 },
        Magic { 0x40404047A0400, 0x2285808020091000, 54, 52224 },
        Magic { 0x8080808760800, 0x400230010010208, 54, 53248 },
        Magic { 0x101010106E1000, 0x542020011482004, 54, 54272 },
        Magic { 0x202020205E2000, 0x808004008200, 54, 55296 },
        Magic { 0x404040403E4000, 0x8900240088251002, 54, 56320 },
        Magic { 0x80808080FE8000, 0x418012000780A104, 52, 57344 },
        Magic { 0x101017F010100, 0x5200400280023020, 52, 61440 },
        Magic { 0x202027C020200, 0xA08A0302002082C0, 54, 65536 },
        Magic { 0x404047A040400, 0x26100280200080, 54, 66560 },
        Magic { 0x8080876080800, 0x3000204200110A00, 54, 67584 },
        Magic { 0x1010106E101000, 0x14080080240180, 54, 68608 },
        Magic { 0x2020205E202000, 0x2000200088410, 54, 69632 },
        Magic { 0x4040403E404000, 0x2802500400421108, 54, 70656 },
        Magic { 0x808080FE808000, 0x80098E100004282, 52, 71680 },
        Magic { 0x1017F01010100, 0xD410400028800094, 52, 75776 },
        Magic { 0x2027C02020200, 0xA800842004804001, 54, 79872 },
        Magic { 0x4047A04040400, 0xD02801000802000, 54, 80896 },
        Magic { 0x8087608080800, 0x3100800800801000, 54, 81920 },
        Magic { 0x10106E10101000, 0x4814012800800480, 54, 82944 },
        Magic { 0x20205E20202000, 0x100801200800400, 54, 83968 },
        Magic { 0x40403E40404000, 0x18211004000802, 54, 84992 },
        Magic { 0x8080FE80808000, 0x102087020000A4, 52, 86016 },
        Magic { 0x17F0101010100, 0x40001044248000, 52, 90112 },
        Magic { 0x27C0202020200, 0x1200050004001, 54, 94208 },
        Magic { 0x47A0404040400, 0x2022200100310042, 54, 95232 },
        Magic { 0x8760808080800, 0x2100181001010020, 54, 96256 },
        Magic { 0x106E1010101000, 0x2002004120008, 54, 97280 },
        Magic { 0x205E2020202000, 0x102001004020008, 54, 98304 },
        Magic { 0x403E4040404000, 0x14048D0020C0001, 54, 99328 },
        Magic { 0x80FE8080808000, 0x1011434004A0001, 52, 100352 },
        Magic { 0x7F010101010100, 0x201422080001500, 52, 104448 },
        Magic { 0x7C020202020200, 0x18C401000A00040, 54, 108544 },
        Magic { 0x7A040404040400, 0xC02210820200, 54, 109568 },
        Magic { 0x76080808080800, 0x21100080180080, 54, 110592 },
        Magic { 0x6E101010101000, 0xB001214280100, 54, 111616 },
        Magic { 0x5E202020202000, 0x8020800200140080, 54, 112640 },
        Magic { 0x3E404040404000, 0x9410800100020080, 54, 113664 },
        Magic { 0xFE808080808000, 0x8000004021000080, 52, 114688 },
        Magic { 0x7E01010101010100, 0x410824108001, 52, 118784 },
        Magic { 0x7E02020202020200, 0x800100880210442, 52, 122880 },
        Magic { 0x7E04040404040400, 0x88060400C191082, 52, 126976 },
        Magic { 0x7E08080808080800, 0x810049810000A21, 52, 131072 },
        Magic { 0x7E10101010101000, 0x2080010A401, 52, 135168 },
        Magic { 0x7E20202020202000, 0x298441000850A, 52, 139264 },
        Magic { 0x7E40404040404000, 0x20809002030144, 52, 143360 },
        Magic { 0x7E80808080808000, 0x2000108044010132, 52, 147456 },
]
pub const rook_table_size = 151552